`timescale 1ns / 1ps


module tb_top;
reg clk;
reg [7:0] a00, a01, a02, a10, a11, a12, a20, a21, a22;
reg [7:0] b00, b01, b02, b10, b11, b12, b20, b21, b22;
wire [7:0] c1,c2,c3,c4,c5,c6,c7,c8,c9;

top uut(
.clk(clk),
.a00(a00), 
.a01(a01), 
.a02(a02), 
.a10(a10), 
.a11(a11), 
.a12(a12), 
.a20(a20), 
.a21(a21), 
.a22(a22),
.b00(b00), 
.b01(b01), 
.b02(b02), 
.b10(b10), 
.b11(b11), 
.b12(b12), 
.b20(b20), 
.b21(b21), 
.b22(b22),
.c1(c1),
.c2(c2),
.c3(c3),
.c4(c4),
.c5(c5),
.c6(c6),
.c7(c7),
.c8(c8),
.c9(c9)
);


initial begin
clk = 0;
a00 = 0;
a01 = 0; 
a02 = 0; 
a10 = 0; 
a11 = 0; 
a12 = 0; 
a20 = 0; 
a21 = 0; 
a22 = 0;
b00 = 0;
b01 = 0; 
b02 = 0; 
b10 = 0; 
b11 = 0; 
b12 = 0; 
b20 = 0; 
b21 = 0; 
b22 = 0;

#50
a00 = 8'b00010000;//0.25
a01 = 8'b10010000; //-0.25
a02 = 8'b00100000; //0.5
a10 = 8'b10100000; //-0.5
a11 = 8'b00110000; //1
a12 = 8'b00110000; //1
a20 = 8'b10111000; //-1.5
a21 = 8'b00111000; //1.5
a22 = 8'b00100111;//0.75
b00 = 8'b10100111;//-0.75
b01 = 8'b00100000; //0.5
b02 = 8'b00110000; //1
b10 = 8'b00110000; //1
b11 = 8'b00010000; //0.25
b12 = 8'b10010000; //-0.25
b20 = 8'b10100000; //-0.5
b21 = 8'b00110000; //1
b22 = 8'b00100000;//0.5

//matrix result should be
//	-0.6875	0.5625	0.5625
//	0.875	1	-0.25
//	2.25	0.375	-1.5

//xa6  x22  x22  
//x2c  x30  x90
//x42  x18  xb8   
end
always
#5 clk = ~clk;
endmodule
